module IU(input wire clk,
			 output wire [7:0] Ins_to_out,
			 output reg [7:0] Operands,
			 input wire  [2:0] enable,
			 output reg[9:0] PC
			);
initial begin
  PC=0;
end
reg [9:0] temp;
reg [7:0] Ins=8'b0;
reg [7:0] ins_mem[1023:0];
initial begin
   ins_mem[0]=8'b11001;
	ins_mem[1]=8'b11111;
	ins_mem[2]=8'b100001;
	ins_mem[3]=8'b1;
	ins_mem[4]=8'b0;
	ins_mem[5]=8'b0;
	ins_mem[6]=8'b100;
	ins_mem[7]=8'b11001;
	ins_mem[8]=8'b100001;
	ins_mem[9]=8'b11001;
	ins_mem[10]=8'b10100;
	ins_mem[11]=8'b101;
	ins_mem[12]=8'b1001;
	ins_mem[13]=8'b11001;
	ins_mem[14]=8'b10111;
	ins_mem[15]=8'b100001;
	ins_mem[16]=8'b10110;
	ins_mem[17]=8'b10100;
	ins_mem[18]=8'b1111;
	ins_mem[19]=8'b11001;
	ins_mem[20]=8'b10111;
	ins_mem[21]=8'b110;
	ins_mem[22]=8'b100001;
	ins_mem[23]=8'b11001;
	ins_mem[24]=8'b10100;
	ins_mem[25]=8'b101;
	ins_mem[26]=8'b1001;
	ins_mem[27]=8'b11001;
	ins_mem[28]=8'b10111;
	ins_mem[29]=8'b10111;
	ins_mem[30]=8'b10111;
	ins_mem[31]=8'b100001;
	ins_mem[32]=8'b10110;
	ins_mem[33]=8'b10100;
	ins_mem[34]=8'b10001;
	ins_mem[35]=8'b11001;
	ins_mem[36]=8'b100;
	ins_mem[37]=8'b11;
	ins_mem[38]=8'b11010000;
	ins_mem[39]=8'b10010001;
	ins_mem[40]=8'b11001;
	ins_mem[41]=8'b10111;
	ins_mem[42]=8'b10111;
	ins_mem[43]=8'b10111;
	ins_mem[44]=8'b1001;
	ins_mem[45]=8'b11;
	ins_mem[46]=8'b11;
	ins_mem[47]=8'b11010000;
	ins_mem[48]=8'b10010001;
	ins_mem[49]=8'b100100;
	ins_mem[50]=8'b10101;
	ins_mem[51]=8'b11100;
	ins_mem[52]=8'b1;
	ins_mem[53]=8'b101011;
	ins_mem[54]=8'b100010;
	ins_mem[55]=8'b10111;
	ins_mem[56]=8'b100;
	ins_mem[57]=8'b11;
	ins_mem[58]=8'b11010000;
	ins_mem[59]=8'b10010001;
	ins_mem[60]=8'b11001;
	ins_mem[61]=8'b10111;
	ins_mem[62]=8'b1010;
	ins_mem[63]=8'b1100;
	ins_mem[64]=8'b11001;
	ins_mem[65]=8'b11111;
	ins_mem[66]=8'b100100;
	ins_mem[67]=8'b100101;
	ins_mem[68]=8'b100001;
	ins_mem[69]=8'b1;
	ins_mem[70]=8'b11;
	ins_mem[71]=8'b11010000;
	ins_mem[72]=8'b10010000;
	ins_mem[73]=8'b11001;
	ins_mem[74]=8'b100001;
	ins_mem[75]=8'b10010;
	ins_mem[76]=8'b10111;
	ins_mem[77]=8'b1001;
	ins_mem[78]=8'b1110;
	ins_mem[79]=8'b11101;
	ins_mem[80]=8'b100001;
	ins_mem[81]=8'b11001;
	ins_mem[82]=8'b100100;
	ins_mem[83]=8'b10000;
	ins_mem[84]=8'b11000;
	ins_mem[85]=8'b1001;
	ins_mem[86]=8'b1011;
	ins_mem[87]=8'b10101;
	ins_mem[88]=8'b11100;
	ins_mem[89]=8'b0;
	ins_mem[90]=8'b11111111;
	ins_mem[91]=8'b1110;
	ins_mem[92]=8'b11000;
	ins_mem[93]=8'b1001;
	ins_mem[94]=8'b1101;
	ins_mem[95]=8'b10101;
	ins_mem[96]=8'b11100;
	ins_mem[97]=8'b0;
	ins_mem[98]=8'b11100010;
	ins_mem[99]=8'b1110;
	ins_mem[100]=8'b1001;
	ins_mem[101]=8'b11001;
	ins_mem[102]=8'b10010;
	ins_mem[103]=8'b11000;
	ins_mem[104]=8'b11110;
	ins_mem[105]=8'b100001;
	ins_mem[106]=8'b11001;
	ins_mem[107]=8'b10100;
	ins_mem[108]=8'b11111;
	ins_mem[109]=8'b11001;
	ins_mem[110]=8'b10010;
	ins_mem[111]=8'b10111;
	ins_mem[112]=8'b100001;
	ins_mem[113]=8'b11001;
	ins_mem[114]=8'b10100;
	ins_mem[115]=8'b110;
	ins_mem[116]=8'b1001;
	ins_mem[117]=8'b100000;
	ins_mem[118]=8'b11101;
	ins_mem[119]=8'b11111;
	ins_mem[120]=8'b11001;
	ins_mem[121]=8'b10010;
	ins_mem[122]=8'b10111;
	ins_mem[123]=8'b100001;
	ins_mem[124]=8'b11001;
	ins_mem[125]=8'b10100;
	ins_mem[126]=8'b1001;
	ins_mem[127]=8'b100000;
	ins_mem[128]=8'b11101;
	ins_mem[129]=8'b11111;
	ins_mem[130]=8'b11001;
	ins_mem[131]=8'b10010;
	ins_mem[132]=8'b1001;
	ins_mem[133]=8'b1110;
	ins_mem[134]=8'b11101;
	ins_mem[135]=8'b100001;
	ins_mem[136]=8'b11001;
	ins_mem[137]=8'b10100;
	ins_mem[138]=8'b110;
	ins_mem[139]=8'b1001;
	ins_mem[140]=8'b100000;
	ins_mem[141]=8'b11101;
	ins_mem[142]=8'b11111;
	ins_mem[143]=8'b11001;
	ins_mem[144]=8'b10010;
	ins_mem[145]=8'b11000;
	ins_mem[146]=8'b100001;
	ins_mem[147]=8'b11001;
	ins_mem[148]=8'b10100;
	ins_mem[149]=8'b110;
	ins_mem[150]=8'b110;
	ins_mem[151]=8'b1001;
	ins_mem[152]=8'b100000;
	ins_mem[153]=8'b11101;
	ins_mem[154]=8'b11111;
	ins_mem[155]=8'b11001;
	ins_mem[156]=8'b10010;
	ins_mem[157]=8'b11000;
	ins_mem[158]=8'b100001;
	ins_mem[159]=8'b11001;
	ins_mem[160]=8'b10100;
	ins_mem[161]=8'b110;
	ins_mem[162]=8'b1001;
	ins_mem[163]=8'b100000;
	ins_mem[164]=8'b11101;
	ins_mem[165]=8'b11111;
	ins_mem[166]=8'b11001;
	ins_mem[167]=8'b10010;
	ins_mem[168]=8'b1001;
	ins_mem[169]=8'b1110;
	ins_mem[170]=8'b11101;
	ins_mem[171]=8'b100001;
	ins_mem[172]=8'b11001;
	ins_mem[173]=8'b10100;
	ins_mem[174]=8'b1001;
	ins_mem[175]=8'b100000;
	ins_mem[176]=8'b11101;
	ins_mem[177]=8'b11111;
	ins_mem[178]=8'b11001;
	ins_mem[179]=8'b10010;
	ins_mem[180]=8'b10111;
	ins_mem[181]=8'b100001;
	ins_mem[182]=8'b11001;
	ins_mem[183]=8'b10100;
	ins_mem[184]=8'b110;
	ins_mem[185]=8'b1001;
	ins_mem[186]=8'b100000;
	ins_mem[187]=8'b11101;
	ins_mem[188]=8'b11111;
	ins_mem[189]=8'b11001;
	ins_mem[190]=8'b10010;
	ins_mem[191]=8'b10111;
	ins_mem[192]=8'b100001;
	ins_mem[193]=8'b11001;
	ins_mem[194]=8'b10100;
	ins_mem[195]=8'b1001;
	ins_mem[196]=8'b100000;
	ins_mem[197]=8'b11101;
	ins_mem[198]=8'b1000;
	ins_mem[199]=8'b1000;
	ins_mem[200]=8'b1000;
	ins_mem[201]=8'b1000;
	ins_mem[202]=8'b11111;
	ins_mem[203]=8'b11001;
	ins_mem[204]=8'b10010;
	ins_mem[205]=8'b100101;
	ins_mem[206]=8'b100010;
	ins_mem[207]=8'b100001;
	ins_mem[208]=8'b10111;
	ins_mem[209]=8'b100100;
	ins_mem[210]=8'b100000;
	ins_mem[211]=8'b10011;
	ins_mem[212]=8'b1110;
	ins_mem[213]=8'b1001;
	ins_mem[214]=8'b11001;
	ins_mem[215]=8'b100011;
	ins_mem[216]=8'b11110;
	ins_mem[217]=8'b10111;
	ins_mem[218]=8'b100001;
	ins_mem[219]=8'b1101;
	ins_mem[220]=8'b10111;
	ins_mem[221]=8'b10111;
	ins_mem[222]=8'b1100;
	ins_mem[223]=8'b11011;
	ins_mem[224]=8'b0;
	ins_mem[225]=8'b1011011;
	ins_mem[226]=8'b11001;
	ins_mem[227]=8'b10111;
	ins_mem[228]=8'b1100;
	ins_mem[229]=8'b1011;
	ins_mem[230]=8'b10111;
	ins_mem[231]=8'b10111;
	ins_mem[232]=8'b1010;
	ins_mem[233]=8'b11001;
	ins_mem[234]=8'b10100;
	ins_mem[235]=8'b1001;
	ins_mem[236]=8'b11001;
	ins_mem[237]=8'b10010;
	ins_mem[238]=8'b100101;
	ins_mem[239]=8'b100010;
	ins_mem[240]=8'b100001;
	ins_mem[241]=8'b10111;
	ins_mem[242]=8'b100100;
	ins_mem[243]=8'b10110;
	ins_mem[244]=8'b10011;
	ins_mem[245]=8'b1110;
	ins_mem[246]=8'b1001;
	ins_mem[247]=8'b100011;
	ins_mem[248]=8'b11101;
	ins_mem[249]=8'b10111;
	ins_mem[250]=8'b10111;
	ins_mem[251]=8'b100001;
	ins_mem[252]=8'b11011;
	ins_mem[253]=8'b0;
	ins_mem[254]=8'b1010011;
	ins_mem[255]=8'b11001;
	ins_mem[256]=8'b10111;
	ins_mem[257]=8'b1100;
	ins_mem[258]=8'b1101;
	ins_mem[259]=8'b1001;
	ins_mem[260]=8'b1110;
	ins_mem[261]=8'b10111;
	ins_mem[262]=8'b11110;
	ins_mem[263]=8'b11100;
	ins_mem[264]=8'b1;
	ins_mem[265]=8'b100010;
	ins_mem[266]=8'b11001;
	ins_mem[267]=8'b10100;
	ins_mem[268]=8'b1001;
	ins_mem[269]=8'b11001;
	ins_mem[270]=8'b10010;
	ins_mem[271]=8'b100101;
	ins_mem[272]=8'b100010;
	ins_mem[273]=8'b100001;
	ins_mem[274]=8'b10111;
	ins_mem[275]=8'b100100;
	ins_mem[276]=8'b10110;
	ins_mem[277]=8'b10011;
	ins_mem[278]=8'b11001;
	ins_mem[279]=8'b100011;
	ins_mem[280]=8'b10111;
	ins_mem[281]=8'b10111;
	ins_mem[282]=8'b100001;
	ins_mem[283]=8'b1101;
	ins_mem[284]=8'b10111;
	ins_mem[285]=8'b10111;
	ins_mem[286]=8'b1100;
	ins_mem[287]=8'b11011;
	ins_mem[288]=8'b1;
	ins_mem[289]=8'b10;
	ins_mem[290]=8'b11001;
	ins_mem[291]=8'b100001;
	ins_mem[292]=8'b10;
	ins_mem[293]=8'b0;
	ins_mem[294]=8'b11110100;
	ins_mem[295]=8'b100100;
	ins_mem[296]=8'b11011;
	ins_mem[297]=8'b0;
	ins_mem[298]=8'b101000;
	ins_mem[299]=8'b100110;
end
assign Ins_to_out=Ins;
always@(negedge clk) begin
	case(enable)
	3'b1: begin
	  Ins=ins_mem[PC];
	  PC<=PC+1;
	end
	3'b10: begin
	  temp=PC;
	  PC[7:0]=ins_mem[temp];
	  temp=temp+1;
	  PC=PC<<8;
	  PC[7:0]<=ins_mem[temp];
	end
	3'b11: begin
	  Operands=ins_mem[PC];
	  PC<=PC+1;
	end
	3'b100:begin
	  PC<=0;
	end
	default: begin
	end
	endcase
end
endmodule
									